module add(a,b,c);
output c;
input a,b;
assign c =a+b;
endmodule
